module block(inp_north, inp_west, clk, rst, outp_south, outp_east, result);
	input [31:0] inp_north, inp_west;
	output reg [31:0] outp_south, outp_east;
	input clk, rst;
	output reg [63:0] result;
	wire [63:0] multi;
	always @(posedge rst or posedge clk) begin
		if(rst) begin
			result <= 0;
			outp_east <= 0;
			outp_south <= 0;
		end
		else begin
			result <= result + multi;
			outp_east <= inp_west;
			outp_south <= inp_north;
		end
	end
	assign multi = inp_north * inp_west;
endmodule

module systolic_array(
	input [31:0] inp_west0, inp_west16, inp_west32, inp_west48, inp_west64, inp_west80, inp_west96, inp_west112,
	             inp_west128, inp_west144, inp_west160, inp_west176, inp_west192, inp_west208, inp_west224, inp_west240,
	input [31:0] inp_north0, inp_north1, inp_north2, inp_north3, inp_north4, inp_north5, inp_north6, inp_north7,
	             inp_north8, inp_north9, inp_north10, inp_north11, inp_north12, inp_north13, inp_north14, inp_north15,
	input clk, rst,
	output reg done,
	output [63:0] result0, result1, result2, result3, result4, result5, result6, result7,
	              result8, result9, result10, result11, result12, result13, result14, result15,
	              result16, result17, result18, result19, result20, result21, result22, result23,
	              result24, result25, result26, result27, result28, result29, result30, result31,
	              result32, result33, result34, result35, result36, result37, result38, result39,
	              result40, result41, result42, result43, result44, result45, result46, result47,
	              result48, result49, result50, result51, result52, result53, result54, result55,
	              result56, result57, result58, result59, result60, result61, result62, result63,
	              result64, result65, result66, result67, result68, result69, result70, result71,
	              result72, result73, result74, result75, result76, result77, result78, result79,
	              result80, result81, result82, result83, result84, result85, result86, result87,
	              result88, result89, result90, result91, result92, result93, result94, result95,
	              result96, result97, result98, result99, result100, result101, result102, result103,
	              result104, result105, result106, result107, result108, result109, result110, result111,
	              result112, result113, result114, result115, result116, result117, result118, result119,
	              result120, result121, result122, result123, result124, result125, result126, result127,
	              result128, result129, result130, result131, result132, result133, result134, result135,
	              result136, result137, result138, result139, result140, result141, result142, result143,
	              result144, result145, result146, result147, result148, result149, result150, result151,
	              result152, result153, result154, result155, result156, result157, result158, result159,
	              result160, result161, result162, result163, result164, result165, result166, result167,
	              result168, result169, result170, result171, result172, result173, result174, result175,
	              result176, result177, result178, result179, result180, result181, result182, result183,
	              result184, result185, result186, result187, result188, result189, result190, result191,
	              result192, result193, result194, result195, result196, result197, result198, result199,
	              result200, result201, result202, result203, result204, result205, result206, result207,
	              result208, result209, result210, result211, result212, result213, result214, result215,
	              result216, result217, result218, result219, result220, result221, result222, result223,
	              result224, result225, result226, result227, result228, result229, result230, result231,
	              result232, result233, result234, result235, result236, result237, result238, result239,
	              result240, result241, result242, result243, result244, result245, result246, result247,
	              result248, result249, result250, result251, result252, result253, result254, result255
);

	// Internal wires
	wire [31:0] outp_south0, outp_south1, outp_south2, outp_south3, outp_south4, outp_south5, outp_south6, outp_south7,
	            outp_south8, outp_south9, outp_south10, outp_south11, outp_south12, outp_south13, outp_south14, outp_south15,
	            outp_south16, outp_south17, outp_south18, outp_south19, outp_south20, outp_south21, outp_south22, outp_south23,
	            outp_south24, outp_south25, outp_south26, outp_south27, outp_south28, outp_south29, outp_south30, outp_south31,
	            outp_south32, outp_south33, outp_south34, outp_south35, outp_south36, outp_south37, outp_south38, outp_south39,
	            outp_south40, outp_south41, outp_south42, outp_south43, outp_south44, outp_south45, outp_south46, outp_south47,
	            outp_south48, outp_south49, outp_south50, outp_south51, outp_south52, outp_south53, outp_south54, outp_south55,
	            outp_south56, outp_south57, outp_south58, outp_south59, outp_south60, outp_south61, outp_south62, outp_south63,
	            outp_south64, outp_south65, outp_south66, outp_south67, outp_south68, outp_south69, outp_south70, outp_south71,
	            outp_south72, outp_south73, outp_south74, outp_south75, outp_south76, outp_south77, outp_south78, outp_south79,
	            outp_south80, outp_south81, outp_south82, outp_south83, outp_south84, outp_south85, outp_south86, outp_south87,
	            outp_south88, outp_south89, outp_south90, outp_south91, outp_south92, outp_south93, outp_south94, outp_south95,
	            outp_south96, outp_south97, outp_south98, outp_south99, outp_south100, outp_south101, outp_south102, outp_south103,
	            outp_south104, outp_south105, outp_south106, outp_south107, outp_south108, outp_south109, outp_south110, outp_south111,
	            outp_south112, outp_south113, outp_south114, outp_south115, outp_south116, outp_south117, outp_south118, outp_south119,
	            outp_south120, outp_south121, outp_south122, outp_south123, outp_south124, outp_south125, outp_south126, outp_south127,
	            outp_south128, outp_south129, outp_south130, outp_south131, outp_south132, outp_south133, outp_south134, outp_south135,
	            outp_south136, outp_south137, outp_south138, outp_south139, outp_south140, outp_south141, outp_south142, outp_south143,
	            outp_south144, outp_south145, outp_south146, outp_south147, outp_south148, outp_south149, outp_south150, outp_south151,
	            outp_south152, outp_south153, outp_south154, outp_south155, outp_south156, outp_south157, outp_south158, outp_south159,
	            outp_south160, outp_south161, outp_south162, outp_south163, outp_south164, outp_south165, outp_south166, outp_south167,
	            outp_south168, outp_south169, outp_south170, outp_south171, outp_south172, outp_south173, outp_south174, outp_south175,
	            outp_south176, outp_south177, outp_south178, outp_south179, outp_south180, outp_south181, outp_south182, outp_south183,
	            outp_south184, outp_south185, outp_south186, outp_south187, outp_south188, outp_south189, outp_south190, outp_south191,
	            outp_south192, outp_south193, outp_south194, outp_south195, outp_south196, outp_south197, outp_south198, outp_south199,
	            outp_south200, outp_south201, outp_south202, outp_south203, outp_south204, outp_south205, outp_south206, outp_south207,
	            outp_south208, outp_south209, outp_south210, outp_south211, outp_south212, outp_south213, outp_south214, outp_south215,
	            outp_south216, outp_south217, outp_south218, outp_south219, outp_south220, outp_south221, outp_south222, outp_south223,
	            outp_south224, outp_south225, outp_south226, outp_south227, outp_south228, outp_south229, outp_south230, outp_south231,
	            outp_south232, outp_south233, outp_south234, outp_south235, outp_south236, outp_south237, outp_south238, outp_south239,
	            outp_south240, outp_south241, outp_south242, outp_south243, outp_south244, outp_south245, outp_south246, outp_south247,
	            outp_south248, outp_south249, outp_south250, outp_south251, outp_south252, outp_south253, outp_south254, outp_south255;

	wire [31:0] outp_east0, outp_east1, outp_east2, outp_east3, outp_east4, outp_east5, outp_east6, outp_east7,
	            outp_east8, outp_east9, outp_east10, outp_east11, outp_east12, outp_east13, outp_east14, outp_east15,
	            outp_east16, outp_east17, outp_east18, outp_east19, outp_east20, outp_east21, outp_east22, outp_east23,
	            outp_east24, outp_east25, outp_east26, outp_east27, outp_east28, outp_east29, outp_east30, outp_east31,
	            outp_east32, outp_east33, outp_east34, outp_east35, outp_east36, outp_east37, outp_east38, outp_east39,
	            outp_east40, outp_east41, outp_east42, outp_east43, outp_east44, outp_east45, outp_east46, outp_east47,
	            outp_east48, outp_east49, outp_east50, outp_east51, outp_east52, outp_east53, outp_east54, outp_east55,
	            outp_east56, outp_east57, outp_east58, outp_east59, outp_east60, outp_east61, outp_east62, outp_east63,
	            outp_east64, outp_east65, outp_east66, outp_east67, outp_east68, outp_east69, outp_east70, outp_east71,
	            outp_east72, outp_east73, outp_east74, outp_east75, outp_east76, outp_east77, outp_east78, outp_east79,
	            outp_east80, outp_east81, outp_east82, outp_east83, outp_east84, outp_east85, outp_east86, outp_east87,
	            outp_east88, outp_east89, outp_east90, outp_east91, outp_east92, outp_east93, outp_east94, outp_east95,
	            outp_east96, outp_east97, outp_east98, outp_east99, outp_east100, outp_east101, outp_east102, outp_east103,
	            outp_east104, outp_east105, outp_east106, outp_east107, outp_east108, outp_east109, outp_east110, outp_east111,
	            outp_east112, outp_east113, outp_east114, outp_east115, outp_east116, outp_east117, outp_east118, outp_east119,
	            outp_east120, outp_east121, outp_east122, outp_east123, outp_east124, outp_east125, outp_east126, outp_east127,
	            outp_east128, outp_east129, outp_east130, outp_east131, outp_east132, outp_east133, outp_east134, outp_east135,
	            outp_east136, outp_east137, outp_east138, outp_east139, outp_east140, outp_east141, outp_east142, outp_east143,
	            outp_east144, outp_east145, outp_east146, outp_east147, outp_east148, outp_east149, outp_east150, outp_east151,
	            outp_east152, outp_east153, outp_east154, outp_east155, outp_east156, outp_east157, outp_east158, outp_east159,
	            outp_east160, outp_east161, outp_east162, outp_east163, outp_east164, outp_east165, outp_east166, outp_east167,
	            outp_east168, outp_east169, outp_east170, outp_east171, outp_east172, outp_east173, outp_east174, outp_east175,
	            outp_east176, outp_east177, outp_east178, outp_east179, outp_east180, outp_east181, outp_east182, outp_east183,
	            outp_east184, outp_east185, outp_east186, outp_east187, outp_east188, outp_east189, outp_east190, outp_east191,
	            outp_east192, outp_east193, outp_east194, outp_east195, outp_east196, outp_east197, outp_east198, outp_east199,
	            outp_east200, outp_east201, outp_east202, outp_east203, outp_east204, outp_east205, outp_east206, outp_east207,
	            outp_east208, outp_east209, outp_east210, outp_east211, outp_east212, outp_east213, outp_east214, outp_east215,
	            outp_east216, outp_east217, outp_east218, outp_east219, outp_east220, outp_east221, outp_east222, outp_east223,
	            outp_east224, outp_east225, outp_east226, outp_east227, outp_east228, outp_east229, outp_east230, outp_east231,
	            outp_east232, outp_east233, outp_east234, outp_east235, outp_east236, outp_east237, outp_east238, outp_east239,
	            outp_east240, outp_east241, outp_east242, outp_east243, outp_east244, outp_east245, outp_east246, outp_east247,
	            outp_east248, outp_east249, outp_east250, outp_east251, outp_east252, outp_east253, outp_east254, outp_east255;

	// Counter for done signal
	reg [6:0] count;

	// Processing Elements (256 PEs for 16x16 array)
	// Row 0
	block P0 (inp_north0, inp_west0, clk, rst, outp_south0, outp_east0, result0);
	block P1 (inp_north1, outp_east0, clk, rst, outp_south1, outp_east1, result1);
	block P2 (inp_north2, outp_east1, clk, rst, outp_south2, outp_east2, result2);
	block P3 (inp_north3, outp_east2, clk, rst, outp_south3, outp_east3, result3);
	block P4 (inp_north4, outp_east3, clk, rst, outp_south4, outp_east4, result4);
	block P5 (inp_north5, outp_east4, clk, rst, outp_south5, outp_east5, result5);
	block P6 (inp_north6, outp_east5, clk, rst, outp_south6, outp_east6, result6);
	block P7 (inp_north7, outp_east6, clk, rst, outp_south7, outp_east7, result7);
	block P8 (inp_north8, outp_east7, clk, rst, outp_south8, outp_east8, result8);
	block P9 (inp_north9, outp_east8, clk, rst, outp_south9, outp_east9, result9);
	block P10 (inp_north10, outp_east9, clk, rst, outp_south10, outp_east10, result10);
	block P11 (inp_north11, outp_east10, clk, rst, outp_south11, outp_east11, result11);
	block P12 (inp_north12, outp_east11, clk, rst, outp_south12, outp_east12, result12);
	block P13 (inp_north13, outp_east12, clk, rst, outp_south13, outp_east13, result13);
	block P14 (inp_north14, outp_east13, clk, rst, outp_south14, outp_east14, result14);
	block P15 (inp_north15, outp_east14, clk, rst, outp_south15, outp_east15, result15);

	// Row 1
	block P16 (outp_south0, inp_west16, clk, rst, outp_south16, outp_east16, result16);
	block P17 (outp_south1, outp_east16, clk, rst, outp_south17, outp_east17, result17);
	block P18 (outp_south2, outp_east17, clk, rst, outp_south18, outp_east18, result18);
	block P19 (outp_south3, outp_east18, clk, rst, outp_south19, outp_east19, result19);
	block P20 (outp_south4, outp_east19, clk, rst, outp_south20, outp_east20, result20);
	block P21 (outp_south5, outp_east20, clk, rst, outp_south21, outp_east21, result21);
	block P22 (outp_south6, outp_east21, clk, rst, outp_south22, outp_east22, result22);
	block P23 (outp_south7, outp_east22, clk, rst, outp_south23, outp_east23, result23);
	block P24 (outp_south8, outp_east23, clk, rst, outp_south24, outp_east24, result24);
	block P25 (outp_south9, outp_east24, clk, rst, outp_south25, outp_east25, result25);
	block P26 (outp_south10, outp_east25, clk, rst, outp_south26, outp_east26, result26);
	block P27 (outp_south11, outp_east26, clk, rst, outp_south27, outp_east27, result27);
	block P28 (outp_south12, outp_east27, clk, rst, outp_south28, outp_east28, result28);
	block P29 (outp_south13, outp_east28, clk, rst, outp_south29, outp_east29, result29);
	block P30 (outp_south14, outp_east29, clk, rst, outp_south30, outp_east30, result30);
	block P31 (outp_south15, outp_east30, clk, rst, outp_south31, outp_east31, result31);

	// Row 2
	block P32 (outp_south16, inp_west32, clk, rst, outp_south32, outp_east32, result32);
	block P33 (outp_south17, outp_east32, clk, rst, outp_south33, outp_east33, result33);
	block P34 (outp_south18, outp_east33, clk, rst, outp_south34, outp_east34, result34);
	block P35 (outp_south19, outp_east34, clk, rst, outp_south35, outp_east35, result35);
	block P36 (outp_south20, outp_east35, clk, rst, outp_south36, outp_east36, result36);
	block P37 (outp_south21, outp_east36, clk, rst, outp_south37, outp_east37, result37);
	block P38 (outp_south22, outp_east37, clk, rst, outp_south38, outp_east38, result38);
	block P39 (outp_south23, outp_east38, clk, rst, outp_south39, outp_east39, result39);
	block P40 (outp_south24, outp_east39, clk, rst, outp_south40, outp_east40, result40);
	block P41 (outp_south25, outp_east40, clk, rst, outp_south41, outp_east41, result41);
	block P42 (outp_south26, outp_east41, clk, rst, outp_south42, outp_east42, result42);
	block P43 (outp_south27, outp_east42, clk, rst, outp_south43, outp_east43, result43);
	block P44 (outp_south28, outp_east43, clk, rst, outp_south44, outp_east44, result44);
	block P45 (outp_south29, outp_east44, clk, rst, outp_south45, outp_east45, result45);
	block P46 (outp_south30, outp_east45, clk, rst, outp_south46, outp_east46, result46);
	block P47 (outp_south31, outp_east46, clk, rst, outp_south47, outp_east47, result47);

	// Row 3
	block P48 (outp_south32, inp_west48, clk, rst, outp_south48, outp_east48, result48);
	block P49 (outp_south33, outp_east48, clk, rst, outp_south49, outp_east49, result49);
	block P50 (outp_south34, outp_east49, clk, rst, outp_south50, outp_east50, result50);
	block P51 (outp_south35, outp_east50, clk, rst, outp_south51, outp_east51, result51);
	block P52 (outp_south36, outp_east51, clk, rst, outp_south52, outp_east52, result52);
	block P53 (outp_south37, outp_east52, clk, rst, outp_south53, outp_east53, result53);
	block P54 (outp_south38, outp_east53, clk, rst, outp_south54, outp_east54, result54);
	block P55 (outp_south39, outp_east54, clk, rst, outp_south55, outp_east55, result55);
	block P56 (outp_south40, outp_east55, clk, rst, outp_south56, outp_east56, result56);
	block P57 (outp_south41, outp_east56, clk, rst, outp_south57, outp_east57, result57);
	block P58 (outp_south42, outp_east57, clk, rst, outp_south58, outp_east58, result58);
	block P59 (outp_south43, outp_east58, clk, rst, outp_south59, outp_east59, result59);
	block P60 (outp_south44, outp_east59, clk, rst, outp_south60, outp_east60, result60);
	block P61 (outp_south45, outp_east60, clk, rst, outp_south61, outp_east61, result61);
	block P62 (outp_south46, outp_east61, clk, rst, outp_south62, outp_east62, result62);
	block P63 (outp_south47, outp_east62, clk, rst, outp_south63, outp_east63, result63);

	// Row 4
	block P64 (outp_south48, inp_west64, clk, rst, outp_south64, outp_east64, result64);
	block P65 (outp_south49, outp_east64, clk, rst, outp_south65, outp_east65, result65);
	block P66 (outp_south50, outp_east65, clk, rst, outp_south66, outp_east66, result66);
	block P67 (outp_south51, outp_east66, clk, rst, outp_south67, outp_east67, result67);
	block P68 (outp_south52, outp_east67, clk, rst, outp_south68, outp_east68, result68);
	block P69 (outp_south53, outp_east68, clk, rst, outp_south69, outp_east69, result69);
	block P70 (outp_south54, outp_east69, clk, rst, outp_south70, outp_east70, result70);
	block P71 (outp_south55, outp_east70, clk, rst, outp_south71, outp_east71, result71);
	block P72 (outp_south56, outp_east71, clk, rst, outp_south72, outp_east72, result72);
	block P73 (outp_south57, outp_east72, clk, rst, outp_south73, outp_east73, result73);
	block P74 (outp_south58, outp_east73, clk, rst, outp_south74, outp_east74, result74);
	block P75 (outp_south59, outp_east74, clk, rst, outp_south75, outp_east75, result75);
	block P76 (outp_south60, outp_east75, clk, rst, outp_south76, outp_east76, result76);
	block P77 (outp_south61, outp_east76, clk, rst, outp_south77, outp_east77, result77);
	block P78 (outp_south62, outp_east77, clk, rst, outp_south78, outp_east78, result78);
	block P79 (outp_south63, outp_east78, clk, rst, outp_south79, outp_east79, result79);

	// Row 5
	block P80 (outp_south64, inp_west80, clk, rst, outp_south80, outp_east80, result80);
	block P81 (outp_south65, outp_east80, clk, rst, outp_south81, outp_east81, result81);
	block P82 (outp_south66, outp_east81, clk, rst, outp_south82, outp_east82, result82);
	block P83 (outp_south67, outp_east82, clk, rst, outp_south83, outp_east83, result83);
	block P84 (outp_south68, outp_east83, clk, rst, outp_south84, outp_east84, result84);
	block P85 (outp_south69, outp_east84, clk, rst, outp_south85, outp_east85, result85);
	block P86 (outp_south70, outp_east85, clk, rst, outp_south86, outp_east86, result86);
	block P87 (outp_south71, outp_east86, clk, rst, outp_south87, outp_east87, result87);
	block P88 (outp_south72, outp_east87, clk, rst, outp_south88, outp_east88, result88);
	block P89 (outp_south73, outp_east88, clk, rst, outp_south89, outp_east89, result89);
	block P90 (outp_south74, outp_east89, clk, rst, outp_south90, outp_east90, result90);
	block P91 (outp_south75, outp_east90, clk, rst, outp_south91, outp_east91, result91);
	block P92 (outp_south76, outp_east91, clk, rst, outp_south92, outp_east92, result92);
	block P93 (outp_south77, outp_east92, clk, rst, outp_south93, outp_east93, result93);
	block P94 (outp_south78, outp_east93, clk, rst, outp_south94, outp_east94, result94);
	block P95 (outp_south79, outp_east94, clk, rst, outp_south95, outp_east95, result95);

	// Row 6
	block P96 (outp_south80, inp_west96, clk, rst, outp_south96, outp_east96, result96);
	block P97 (outp_south81, outp_east96, clk, rst, outp_south97, outp_east97, result97);
	block P98 (outp_south82, outp_east97, clk, rst, outp_south98, outp_east98, result98);
	block P99 (outp_south83, outp_east98, clk, rst, outp_south99, outp_east99, result99);
	block P100 (outp_south84, outp_east99, clk, rst, outp_south100, outp_east100, result100);
	block P101 (outp_south85, outp_east100, clk, rst, outp_south101, outp_east101, result101);
	block P102 (outp_south86, outp_east101, clk, rst, outp_south102, outp_east102, result102);
	block P103 (outp_south87, outp_east102, clk, rst, outp_south103, outp_east103, result103);
	block P104 (outp_south88, outp_east103, clk, rst, outp_south104, outp_east104, result104);
	block P105 (outp_south89, outp_east104, clk, rst, outp_south105, outp_east105, result105);
	block P106 (outp_south90, outp_east105, clk, rst, outp_south106, outp_east106, result106);
	block P107 (outp_south91, outp_east106, clk, rst, outp_south107, outp_east107, result107);
	block P108 (outp_south92, outp_east107, clk, rst, outp_south108, outp_east108, result108);
	block P109 (outp_south93, outp_east108, clk, rst, outp_south109, outp_east109, result109);
	block P110 (outp_south94, outp_east109, clk, rst, outp_south110, outp_east110, result110);
	block P111 (outp_south95, outp_east110, clk, rst, outp_south111, outp_east111, result111);

	// Row 7
	block P112 (outp_south96, inp_west112, clk, rst, outp_south112, outp_east112, result112);
	block P113 (outp_south97, outp_east112, clk, rst, outp_south113, outp_east113, result113);
	block P114 (outp_south98, outp_east113, clk, rst, outp_south114, outp_east114, result114);
	block P115 (outp_south99, outp_east114, clk, rst, outp_south115, outp_east115, result115);
	block P116 (outp_south100, outp_east115, clk, rst, outp_south116, outp_east116, result116);
	block P117 (outp_south101, outp_east116, clk, rst, outp_south117, outp_east117, result117);
	block P118 (outp_south102, outp_east117, clk, rst, outp_south118, outp_east118, result118);
	block P119 (outp_south103, outp_east118, clk, rst, outp_south119, outp_east119, result119);
	block P120 (outp_south104, outp_east119, clk, rst, outp_south120, outp_east120, result120);
	block P121 (outp_south105, outp_east120, clk, rst, outp_south121, outp_east121, result121);
	block P122 (outp_south106, outp_east121, clk, rst, outp_south122, outp_east122, result122);
	block P123 (outp_south107, outp_east122, clk, rst, outp_south123, outp_east123, result123);
	block P124 (outp_south108, outp_east123, clk, rst, outp_south124, outp_east124, result124);
	block P125 (outp_south109, outp_east124, clk, rst, outp_south125, outp_east125, result125);
	block P126 (outp_south110, outp_east125, clk, rst, outp_south126, outp_east126, result126);
	block P127 (outp_south111, outp_east126, clk, rst, outp_south127, outp_east127, result127);

	// Row 8
	block P128 (outp_south112, inp_west128, clk, rst, outp_south128, outp_east128, result128);
	block P129 (outp_south113, outp_east128, clk, rst, outp_south129, outp_east129, result129);
	block P130 (outp_south114, outp_east129, clk, rst, outp_south130, outp_east130, result130);
	block P131 (outp_south115, outp_east130, clk, rst, outp_south131, outp_east131, result131);
	block P132 (outp_south116, outp_east131, clk, rst, outp_south132, outp_east132, result132);
	block P133 (outp_south117, outp_east132, clk, rst, outp_south133, outp_east133, result133);
	block P134 (outp_south118, outp_east133, clk, rst, outp_south134, outp_east134, result134);
	block P135 (outp_south119, outp_east134, clk, rst, outp_south135, outp_east135, result135);
	block P136 (outp_south120, outp_east135, clk, rst, outp_south136, outp_east136, result136);
	block P137 (outp_south121, outp_east136, clk, rst, outp_south137, outp_east137, result137);
	block P138 (outp_south122, outp_east137, clk, rst, outp_south138, outp_east138, result138);
	block P139 (outp_south123, outp_east138, clk, rst, outp_south139, outp_east139, result139);
	block P140 (outp_south124, outp_east139, clk, rst, outp_south140, outp_east140, result140);
	block P141 (outp_south125, outp_east140, clk, rst, outp_south141, outp_east141, result141);
	block P142 (outp_south126, outp_east141, clk, rst, outp_south142, outp_east142, result142);
	block P143 (outp_south127, outp_east142, clk, rst, outp_south143, outp_east143, result143);

	// Row 9
	block P144 (outp_south128, inp_west144, clk, rst, outp_south144, outp_east144, result144);
	block P145 (outp_south129, outp_east144, clk, rst, outp_south145, outp_east145, result145);
	block P146 (outp_south130, outp_east145, clk, rst, outp_south146, outp_east146, result146);
	block P147 (outp_south131, outp_east146, clk, rst, outp_south147, outp_east147, result147);
	block P148 (outp_south132, outp_east147, clk, rst, outp_south148, outp_east148, result148);
	block P149 (outp_south133, outp_east148, clk, rst, outp_south149, outp_east149, result149);
	block P150 (outp_south134, outp_east149, clk, rst, outp_south150, outp_east150, result150);
	block P151 (outp_south135, outp_east150, clk, rst, outp_south151, outp_east151, result151);
	block P152 (outp_south136, outp_east151, clk, rst, outp_south152, outp_east152, result152);
	block P153 (outp_south137, outp_east152, clk, rst, outp_south153, outp_east153, result153);
	block P154 (outp_south138, outp_east153, clk, rst, outp_south154, outp_east154, result154);
	block P155 (outp_south139, outp_east154, clk, rst, outp_south155, outp_east155, result155);
	block P156 (outp_south140, outp_east155, clk, rst, outp_south156, outp_east156, result156);
	block P157 (outp_south141, outp_east156, clk, rst, outp_south157, outp_east157, result157);
	block P158 (outp_south142, outp_east157, clk, rst, outp_south158, outp_east158, result158);
	block P159 (outp_south143, outp_east158, clk, rst, outp_south159, outp_east159, result159);

	// Row 10
	block P160 (outp_south144, inp_west160, clk, rst, outp_south160, outp_east160, result160);
	block P161 (outp_south145, outp_east160, clk, rst, outp_south161, outp_east161, result161);
	block P162 (outp_south146, outp_east161, clk, rst, outp_south162, outp_east162, result162);
	block P163 (outp_south147, outp_east162, clk, rst, outp_south163, outp_east163, result163);
	block P164 (outp_south148, outp_east163, clk, rst, outp_south164, outp_east164, result164);
	block P165 (outp_south149, outp_east164, clk, rst, outp_south165, outp_east165, result165);
	block P166 (outp_south150, outp_east165, clk, rst, outp_south166, outp_east166, result166);
	block P167 (outp_south151, outp_east166, clk, rst, outp_south167, outp_east167, result167);
	block P168 (outp_south152, outp_east167, clk, rst, outp_south168, outp_east168, result168);
	block P169 (outp_south153, outp_east168, clk, rst, outp_south169, outp_east169, result169);
	block P170 (outp_south154, outp_east169, clk, rst, outp_south170, outp_east170, result170);
	block P171 (outp_south155, outp_east170, clk, rst, outp_south171, outp_east171, result171);
	block P172 (outp_south156, outp_east171, clk, rst, outp_south172, outp_east172, result172);
	block P173 (outp_south157, outp_east172, clk, rst, outp_south173, outp_east173, result173);
	block P174 (outp_south158, outp_east173, clk, rst, outp_south174, outp_east174, result174);
	block P175 (outp_south159, outp_east174, clk, rst, outp_south175, outp_east175, result175);

	// Row 11
	block P176 (outp_south160, inp_west176, clk, rst, outp_south176, outp_east176, result176);
	block P177 (outp_south161, outp_east176, clk, rst, outp_south177, outp_east177, result177);
	block P178 (outp_south162, outp_east177, clk, rst, outp_south178, outp_east178, result178);
	block P179 (outp_south163, outp_east178, clk, rst, outp_south179, outp_east179, result179);
	block P180 (outp_south164, outp_east179, clk, rst, outp_south180, outp_east180, result180);
	block P181 (outp_south165, outp_east180, clk, rst, outp_south181, outp_east181, result181);
	block P182 (outp_south166, outp_east181, clk, rst, outp_south182, outp_east182, result182);
	block P183 (outp_south167, outp_east182, clk, rst, outp_south183, outp_east183, result183);
	block P184 (outp_south168, outp_east183, clk, rst, outp_south184, outp_east184, result184);
	block P185 (outp_south169, outp_east184, clk, rst, outp_south185, outp_east185, result185);
	block P186 (outp_south170, outp_east185, clk, rst, outp_south186, outp_east186, result186);
	block P187 (outp_south171, outp_east186, clk, rst, outp_south187, outp_east187, result187);
	block P188 (outp_south172, outp_east187, clk, rst, outp_south188, outp_east188, result188);
	block P189 (outp_south173, outp_east188, clk, rst, outp_south189, outp_east189, result189);
	block P190 (outp_south174, outp_east189, clk, rst, outp_south190, outp_east190, result190);
	block P191 (outp_south175, outp_east190, clk, rst, outp_south191, outp_east191, result191);

	// Row 12
	block P192 (outp_south176, inp_west192, clk, rst, outp_south192, outp_east192, result192);
	block P193 (outp_south177, outp_east192, clk, rst, outp_south193, outp_east193, result193);
	block P194 (outp_south178, outp_east193, clk, rst, outp_south194, outp_east194, result194);
	block P195 (outp_south179, outp_east194, clk, rst, outp_south195, outp_east195, result195);
	block P196 (outp_south180, outp_east195, clk, rst, outp_south196, outp_east196, result196);
	block P197 (outp_south181, outp_east196, clk, rst, outp_south197, outp_east197, result197);
	block P198 (outp_south182, outp_east197, clk, rst, outp_south198, outp_east198, result198);
	block P199 (outp_south183, outp_east198, clk, rst, outp_south199, outp_east199, result199);
	block P200 (outp_south184, outp_east199, clk, rst, outp_south200, outp_east200, result200);
	block P201 (outp_south185, outp_east200, clk, rst, outp_south201, outp_east201, result201);
	block P202 (outp_south186, outp_east201, clk, rst, outp_south202, outp_east202, result202);
	block P203 (outp_south187, outp_east202, clk, rst, outp_south203, outp_east203, result203);
	block P204 (outp_south188, outp_east203, clk, rst, outp_south204, outp_east204, result204);
	block P205 (outp_south189, outp_east204, clk, rst, outp_south205, outp_east205, result205);
	block P206 (outp_south190, outp_east205, clk, rst, outp_south206, outp_east206, result206);
	block P207 (outp_south191, outp_east206, clk, rst, outp_south207, outp_east207, result207);

	// Row 13
	block P208 (outp_south192, inp_west208, clk, rst, outp_south208, outp_east208, result208);
	block P209 (outp_south193, outp_east208, clk, rst, outp_south209, outp_east209, result209);
	block P210 (outp_south194, outp_east209, clk, rst, outp_south210, outp_east210, result210);
	block P211 (outp_south195, outp_east210, clk, rst, outp_south211, outp_east211, result211);
	block P212 (outp_south196, outp_east211, clk, rst, outp_south212, outp_east212, result212);
	block P213 (outp_south197, outp_east212, clk, rst, outp_south213, outp_east213, result213);
	block P214 (outp_south198, outp_east213, clk, rst, outp_south214, outp_east214, result214);
	block P215 (outp_south199, outp_east214, clk, rst, outp_south215, outp_east215, result215);
	block P216 (outp_south200, outp_east215, clk, rst, outp_south216, outp_east216, result216);
	block P217 (outp_south201, outp_east216, clk, rst, outp_south217, outp_east217, result217);
	block P218 (outp_south202, outp_east217, clk, rst, outp_south218, outp_east218, result218);
	block P219 (outp_south203, outp_east218, clk, rst, outp_south219, outp_east219, result219);
	block P220 (outp_south204, outp_east219, clk, rst, outp_south220, outp_east220, result220);
	block P221 (outp_south205, outp_east220, clk, rst, outp_south221, outp_east221, result221);
	block P222 (outp_south206, outp_east221, clk, rst, outp_south222, outp_east222, result222);
	block P223 (outp_south207, outp_east222, clk, rst, outp_south223, outp_east223, result223);

	// Row 14
	block P224 (outp_south208, inp_west224, clk, rst, outp_south224, outp_east224, result224);
	block P225 (outp_south209, outp_east224, clk, rst, outp_south225, outp_east225, result225);
	block P226 (outp_south210, outp_east225, clk, rst, outp_south226, outp_east226, result226);
	block P227 (outp_south211, outp_east226, clk, rst, outp_south227, outp_east227, result227);
	block P228 (outp_south212, outp_east227, clk, rst, outp_south228, outp_east228, result228);
	block P229 (outp_south213, outp_east228, clk, rst, outp_south229, outp_east229, result229);
	block P230 (outp_south214, outp_east229, clk, rst, outp_south230, outp_east230, result230);
	block P231 (outp_south215, outp_east230, clk, rst, outp_south231, outp_east231, result231);
	block P232 (outp_south216, outp_east231, clk, rst, outp_south232, outp_east232, result232);
	block P233 (outp_south217, outp_east232, clk, rst, outp_south233, outp_east233, result233);
	block P234 (outp_south218, outp_east233, clk, rst, outp_south234, outp_east234, result234);
	block P235 (outp_south219, outp_east234, clk, rst, outp_south235, outp_east235, result235);
	block P236 (outp_south220, outp_east235, clk, rst, outp_south236, outp_east236, result236);
	block P237 (outp_south221, outp_east236, clk, rst, outp_south237, outp_east237, result237);
	block P238 (outp_south222, outp_east237, clk, rst, outp_south238, outp_east238, result238);
	block P239 (outp_south223, outp_east238, clk, rst, outp_south239, outp_east239, result239);

	// Row 15
	block P240 (outp_south224, inp_west240, clk, rst, outp_south240, outp_east240, result240);
	block P241 (outp_south225, outp_east240, clk, rst, outp_south241, outp_east241, result241);
	block P242 (outp_south226, outp_east241, clk, rst, outp_south242, outp_east242, result242);
	block P243 (outp_south227, outp_east242, clk, rst, outp_south243, outp_east243, result243);
	block P244 (outp_south228, outp_east243, clk, rst, outp_south244, outp_east244, result244);
	block P245 (outp_south229, outp_east244, clk, rst, outp_south245, outp_east245, result245);
	block P246 (outp_south230, outp_east245, clk, rst, outp_south246, outp_east246, result246);
	block P247 (outp_south231, outp_east246, clk, rst, outp_south247, outp_east247, result247);
	block P248 (outp_south232, outp_east247, clk, rst, outp_south248, outp_east248, result248);
	block P249 (outp_south233, outp_east248, clk, rst, outp_south249, outp_east249, result249);
	block P250 (outp_south234, outp_east249, clk, rst, outp_south250, outp_east250, result250);
	block P251 (outp_south235, outp_east250, clk, rst, outp_south251, outp_east251, result251);
	block P252 (outp_south236, outp_east251, clk, rst, outp_south252, outp_east252, result252);
	block P253 (outp_south237, outp_east252, clk, rst, outp_south253, outp_east253, result253);
	block P254 (outp_south238, outp_east253, clk, rst, outp_south254, outp_east254, result254);
	block P255 (outp_south239, outp_east254, clk, rst, outp_south255, outp_east255, result255);

	// Done signal logic
	always @(posedge clk or posedge rst) begin
		if(rst) begin
			done <= 0;
			count <= 0;
		end
		else begin
			if(count == 46) begin
				done <= 1;
				count <= 0;
			end
			else begin
				done <= 0;
				count <= count + 1;
			end
		end
	end

endmodule
